../register_space.vh