 module ADC_Deserializer(  input wire reset,  input wire data_a,  input wire data_b,  input wire data_c,  input wire data_d,  input wire data_clk,  input wire frame_clk,  output reg [9:0] deser_a,  output reg [9:0] deser_b,  output reg [9:0] deser_c,  output reg [9:0] deser_d);wire q_a, q_b, q_c, q_d;always @(posedge frame_clk)begin  deser_a <= q_a;  deser_b <= q_b;  deser_c <= q_c;  deser_d <= q_d;endADC_ShiftRegister channel_A_ShiftRegister (  .aclr ( reset ),  .clock ( data_clk ),  .shiftin ( data_a ),  .q ( q_a )  );ADC_ShiftRegister channel_B_ShiftRegister (  .aclr ( reset ),  .clock ( data_clk ),  .shiftin ( data_b ),  .q ( q_b )  );ADC_ShiftRegister channel_C_ShiftRegister (  .aclr ( reset ),  .clock ( data_clk ),  .shiftin ( data_c ),  .q ( q_c )  );ADC_ShiftRegister channel_D_ShiftRegister (  .aclr ( reset ),  .clock ( data_clk ),  .shiftin ( data_d ),  .q ( q_d )  );endmodule