`timescale 1 ns / 1 psmodule switch_debounce(  input clk,  input switch_in,  output wire switch_out);assign switch_out = (((fast_enable && fast_out) || hit1) && jitter_filter);reg jitter_filter;reg [10:0]jitter_counter;reg switch_prev;always @(posedge clk) begin  switch_prev <= switch_in;  if (switch_prev != switch_in)    jitter_counter <= 0;  else if (jitter_counter == 11'hFFFFF)    jitter_filter <= switch_in;  else    jitter_counter <= jitter_counter + 1;endreg hit1;reg fast_enable;reg [25:0]cnt;always @(posedge clk) begin  if (jitter_filter == 1) begin    if (cnt == 0) begin      hit1 <= 1;      cnt <= 1;    end    else if (cnt == 26'hFFFFFFF) begin      fast_enable <= 1;      hit1 <= 0;    end    else begin      fast_enable <= 0;      cnt <= cnt + 1;      hit1 <= 0;    end  end  else begin    fast_enable <= 0;    cnt = 0;    hit1 <= 0;  endendreg [24:0]fast_cycle;reg fast_out;always @(posedge clk)begin  fast_cycle <= fast_cycle + 1;  if (fast_cycle == 25'hFFFFFFF)    fast_out <= 1;  else    fast_out <= 0;endendmodule