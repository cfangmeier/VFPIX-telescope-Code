../instruction_set.vh