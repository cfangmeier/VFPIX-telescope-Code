`timescale 1 ns / 1 ps

module seven_segment_display
(
  input clk,
  input [15:0]num_in,
  output reg [6:0]hex0,
  output reg [6:0]hex1,
  output reg [6:0]hex2,
  output reg [6:0]hex3
);

//digit format
//dig[0] : A, top
//dig[1] : B, top/right
//dig[2] : C, bottom/right
//dig[3] : D, bottom
//dig[4] : E, bottom/left
//dig[5] : F, top/left
//dig[6] : G, middle

always @(posedge clk) begin
  case(num_in[3:0])
    4'b0000: hex0 = 7'b1000000; //0
    4'b0001: hex0 = 7'b1111001; //1
    4'b0010: hex0 = 7'b0100100; //2
    4'b0011: hex0 = 7'b0110000; //3
    4'b0100: hex0 = 7'b0011001; //4
    4'b0101: hex0 = 7'b0010010; //5
    4'b0110: hex0 = 7'b0000010; //6
    4'b0111: hex0 = 7'b1111000; //7
    4'b1000: hex0 = 7'b0000000; //8
    4'b1001: hex0 = 7'b0010000; //9
    4'b1010: hex0 = 7'b0001000; //A
    4'b1011: hex0 = 7'b0000011; //b
    4'b1100: hex0 = 7'b1000110; //C
    4'b1101: hex0 = 7'b0100001; //d
    4'b1110: hex0 = 7'b0000110; //E
    4'b1111: hex0 = 7'b0001110; //F
  endcase
  case(num_in[7:4])
    4'b0000: hex1 = 7'b1000000; //0
    4'b0001: hex1 = 7'b1111001; //1
    4'b0010: hex1 = 7'b0100100; //2
    4'b0011: hex1 = 7'b0110000; //3
    4'b0100: hex1 = 7'b0011001; //4
    4'b0101: hex1 = 7'b0010010; //5
    4'b0110: hex1 = 7'b0000010; //6
    4'b0111: hex1 = 7'b1111000; //7
    4'b1000: hex1 = 7'b0000000; //8
    4'b1001: hex1 = 7'b0010000; //9
    4'b1010: hex1 = 7'b0001000; //A
    4'b1011: hex1 = 7'b0000011; //b
    4'b1100: hex1 = 7'b1000110; //C
    4'b1101: hex1 = 7'b0100001; //d
    4'b1110: hex1 = 7'b0000110; //E
    4'b1111: hex1 = 7'b0001110; //F
  endcase
  case(num_in[11:8])
    4'b0000: hex2 = 7'b1000000; //0
    4'b0001: hex2 = 7'b1111001; //1
    4'b0010: hex2 = 7'b0100100; //2
    4'b0011: hex2 = 7'b0110000; //3
    4'b0100: hex2 = 7'b0011001; //4
    4'b0101: hex2 = 7'b0010010; //5
    4'b0110: hex2 = 7'b0000010; //6
    4'b0111: hex2 = 7'b1111000; //7
    4'b1000: hex2 = 7'b0000000; //8
    4'b1001: hex2 = 7'b0010000; //9
    4'b1010: hex2 = 7'b0001000; //A
    4'b1011: hex2 = 7'b0000011; //b
    4'b1100: hex2 = 7'b1000110; //C
    4'b1101: hex2 = 7'b0100001; //d
    4'b1110: hex2 = 7'b0000110; //E
    4'b1111: hex2 = 7'b0001110; //F
  endcase
  case(num_in[15:12])
    4'b0000: hex3 = 7'b1000000; //0
    4'b0001: hex3 = 7'b1111001; //1
    4'b0010: hex3 = 7'b0100100; //2
    4'b0011: hex3 = 7'b0110000; //3
    4'b0100: hex3 = 7'b0011001; //4
    4'b0101: hex3 = 7'b0010010; //5
    4'b0110: hex3 = 7'b0000010; //6
    4'b0111: hex3 = 7'b1111000; //7
    4'b1000: hex3 = 7'b0000000; //8
    4'b1001: hex3 = 7'b0010000; //9
    4'b1010: hex3 = 7'b0001000; //A
    4'b1011: hex3 = 7'b0000011; //b
    4'b1100: hex3 = 7'b1000110; //C
    4'b1101: hex3 = 7'b0100001; //d
    4'b1110: hex3 = 7'b0000110; //E
    4'b1111: hex3 = 7'b0001110; //F
  endcase
end

endmodule
